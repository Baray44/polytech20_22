// my_ISSP.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module my_ISSP (
		input  wire       source_clk, // source_clk.clk
		output wire [8:0] source      //    sources.source
	);

	altsource_probe_top #(
		.sld_auto_instance_index ("YES"),
		.sld_instance_index      (0),
		.instance_id             ("my"),
		.probe_width             (0),
		.source_width            (9),
		.source_initial_value    ("0"),
		.enable_metastability    ("YES")
	) in_system_sources_probes_0 (
		.source     (source),     //    sources.source
		.source_clk (source_clk), // source_clk.clk
		.source_ena (1'b1)        // (terminated)
	);

endmodule
