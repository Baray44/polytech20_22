// Lab4_sys.v

// Generated using ACDS version 16.1 203

`timescale 1 ps / 1 ps
module Lab4_sys (
		input  wire       clk_clk,          //       clk.clk
		output wire [7:0] d_slave_export,   //   d_slave.export
		input  wire [7:0] data_d_export,    //    data_d.export
		output wire [7:0] dd_slave_export,  //  dd_slave.export
		output wire [7:0] def_slave_export, // def_slave.export
		input  wire       reset_reset_n     //     reset.reset_n
	);

	wire        my_master_0_m0_waitrequest;                   // mm_interconnect_0:my_master_0_m0_waitrequest -> my_master_0:avm_m0_waitrequest
	wire  [7:0] my_master_0_m0_address;                       // my_master_0:avm_m0_address -> mm_interconnect_0:my_master_0_m0_address
	wire        my_master_0_m0_write;                         // my_master_0:avm_m0_write -> mm_interconnect_0:my_master_0_m0_write
	wire  [7:0] my_master_0_m0_writedata;                     // my_master_0:avm_m0_writedata -> mm_interconnect_0:my_master_0_m0_writedata
	wire        mm_interconnect_0_my_slave_0_s0_waitrequest;  // my_slave_0:avs_s0_waitrequest -> mm_interconnect_0:my_slave_0_s0_waitrequest
	wire        mm_interconnect_0_my_slave_0_s0_write;        // mm_interconnect_0:my_slave_0_s0_write -> my_slave_0:avs_s0_write
	wire  [7:0] mm_interconnect_0_my_slave_0_s0_writedata;    // mm_interconnect_0:my_slave_0_s0_writedata -> my_slave_0:avs_s0_writedata
	wire        mm_interconnect_0_my_slave_1_s0_waitrequest;  // my_slave_1:avs_s0_waitrequest -> mm_interconnect_0:my_slave_1_s0_waitrequest
	wire        mm_interconnect_0_my_slave_1_s0_write;        // mm_interconnect_0:my_slave_1_s0_write -> my_slave_1:avs_s0_write
	wire  [7:0] mm_interconnect_0_my_slave_1_s0_writedata;    // mm_interconnect_0:my_slave_1_s0_writedata -> my_slave_1:avs_s0_writedata
	wire        mm_interconnect_0_my_dslave_0_s0_waitrequest; // my_Dslave_0:avs_s0_waitrequest -> mm_interconnect_0:my_Dslave_0_s0_waitrequest
	wire        mm_interconnect_0_my_dslave_0_s0_write;       // mm_interconnect_0:my_Dslave_0_s0_write -> my_Dslave_0:avs_s0_write
	wire  [7:0] mm_interconnect_0_my_dslave_0_s0_writedata;   // mm_interconnect_0:my_Dslave_0_s0_writedata -> my_Dslave_0:avs_s0_writedata

	my_Dslave my_dslave_0 (
		.csi_clk            (clk_clk),                                      //         clock.clk
		.rsi_reset          (~reset_reset_n),                               //         reset.reset
		.avs_s0_writedata   (mm_interconnect_0_my_dslave_0_s0_writedata),   //            s0.writedata
		.avs_s0_write       (mm_interconnect_0_my_dslave_0_s0_write),       //              .write
		.avs_s0_waitrequest (mm_interconnect_0_my_dslave_0_s0_waitrequest), //              .waitrequest
		.coe_s0_Dout        (def_slave_export)                              // conduit_end_0.export
	);

	my_master my_master_0 (
		.csi_clk            (clk_clk),                    //         clock.clk
		.rsi_reset          (~reset_reset_n),             //         reset.reset
		.avm_m0_address     (my_master_0_m0_address),     //            m0.address
		.avm_m0_write       (my_master_0_m0_write),       //              .write
		.avm_m0_writedata   (my_master_0_m0_writedata),   //              .writedata
		.avm_m0_waitrequest (my_master_0_m0_waitrequest), //              .waitrequest
		.coe_c0_DA          (data_d_export)               // conduit_end_0.export
	);

	my_slave my_slave_0 (
		.csi_clk            (clk_clk),                                     //         clock.clk
		.rsi_reset          (~reset_reset_n),                              //         reset.reset
		.avs_s0_writedata   (mm_interconnect_0_my_slave_0_s0_writedata),   //            s0.writedata
		.avs_s0_write       (mm_interconnect_0_my_slave_0_s0_write),       //              .write
		.avs_s0_waitrequest (mm_interconnect_0_my_slave_0_s0_waitrequest), //              .waitrequest
		.coe_s0_Dout        (d_slave_export)                               // conduit_end_0.export
	);

	my_slave my_slave_1 (
		.csi_clk            (clk_clk),                                     //         clock.clk
		.rsi_reset          (~reset_reset_n),                              //         reset.reset
		.avs_s0_writedata   (mm_interconnect_0_my_slave_1_s0_writedata),   //            s0.writedata
		.avs_s0_write       (mm_interconnect_0_my_slave_1_s0_write),       //              .write
		.avs_s0_waitrequest (mm_interconnect_0_my_slave_1_s0_waitrequest), //              .waitrequest
		.coe_s0_Dout        (dd_slave_export)                              // conduit_end_0.export
	);

	Lab4_sys_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                      //                               clk_0_clk.clk
		.my_master_0_reset_reset_bridge_in_reset_reset (~reset_reset_n),                               // my_master_0_reset_reset_bridge_in_reset.reset
		.my_master_0_m0_address                        (my_master_0_m0_address),                       //                          my_master_0_m0.address
		.my_master_0_m0_waitrequest                    (my_master_0_m0_waitrequest),                   //                                        .waitrequest
		.my_master_0_m0_write                          (my_master_0_m0_write),                         //                                        .write
		.my_master_0_m0_writedata                      (my_master_0_m0_writedata),                     //                                        .writedata
		.my_Dslave_0_s0_write                          (mm_interconnect_0_my_dslave_0_s0_write),       //                          my_Dslave_0_s0.write
		.my_Dslave_0_s0_writedata                      (mm_interconnect_0_my_dslave_0_s0_writedata),   //                                        .writedata
		.my_Dslave_0_s0_waitrequest                    (mm_interconnect_0_my_dslave_0_s0_waitrequest), //                                        .waitrequest
		.my_slave_0_s0_write                           (mm_interconnect_0_my_slave_0_s0_write),        //                           my_slave_0_s0.write
		.my_slave_0_s0_writedata                       (mm_interconnect_0_my_slave_0_s0_writedata),    //                                        .writedata
		.my_slave_0_s0_waitrequest                     (mm_interconnect_0_my_slave_0_s0_waitrequest),  //                                        .waitrequest
		.my_slave_1_s0_write                           (mm_interconnect_0_my_slave_1_s0_write),        //                           my_slave_1_s0.write
		.my_slave_1_s0_writedata                       (mm_interconnect_0_my_slave_1_s0_writedata),    //                                        .writedata
		.my_slave_1_s0_waitrequest                     (mm_interconnect_0_my_slave_1_s0_waitrequest)   //                                        .waitrequest
	);

endmodule
